ntm_addressing_content.vhd
ntm_addressing_location.vhd
ntm_convolution.vhd
ntm_interpolation.vhd
ntm_reading.vhd
ntm_sharpening.vhd
ntm_writing.vhd