// File vhdl/dnc/write_heads/dnc_write_vector.vhd translated with vhd2vl v2.5 VHDL to Verilog RTL translator
// vhd2vl settings:
//  * Verilog Module Declaration Style: 1995

// vhd2vl is Free (libre) Software:
//   Copyright (C) 2001 Vincenzo Liguori - Ocean Logic Pty Ltd
//     http://www.ocean-logic.com
//   Modifications Copyright (C) 2006 Mark Gonzales - PMC Sierra Inc
//   Modifications (C) 2010 Shankar Giri
//   Modifications Copyright (C) 2002, 2005, 2008-2010, 2015 Larry Doolittle - LBNL
//     http://doolittle.icarus.com/~larry/vhd2vl/
//
//   vhd2vl comes with ABSOLUTELY NO WARRANTY.  Always check the resulting
//   Verilog for correctness, ideally with a formal verification tool.
//
//   You are welcome to redistribute vhd2vl under certain conditions.
//   See the license (GPLv2) file included with the source for details.

// The result of translation follows.  Its copyright status should be
// considered unchanged from the original VHDL.

//------------------------------------------------------------------------------
//                                            __ _      _     _               --
//                                           / _(_)    | |   | |              --
//                __ _ _   _  ___  ___ _ __ | |_ _  ___| | __| |              --
//               / _` | | | |/ _ \/ _ \ '_ \|  _| |/ _ \ |/ _` |              --
//              | (_| | |_| |  __/  __/ | | | | | |  __/ | (_| |              --
//               \__, |\__,_|\___|\___|_| |_|_| |_|\___|_|\__,_|              --
//                  | |                                                       --
//                  |_|                                                       --
//                                                                            --
//                                                                            --
//              Peripheral-NTM for MPSoC                                      --
//              Neural Turing Machine for MPSoC                               --
//                                                                            --
//------------------------------------------------------------------------------
// Copyright (c) 2020-2021 by the author(s)
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
//------------------------------------------------------------------------------
// Author(s):
//   Paco Reina Campo <pacoreinacampo@queenfield.tech>
// no timescale needed

module dnc_write_vector(
CLK,
RST,
START,
READY,
V_IN_ENABLE,
V_OUT_ENABLE,
SIZE_W_IN,
V_IN,
V_OUT
);

parameter [31:0] DATA_SIZE=512;
// GLOBAL
input CLK;
input RST;
// CONTROL
input START;
output READY;
input V_IN_ENABLE;
// for k in 0 to W-1
output V_OUT_ENABLE;
// for k in 0 to W-1
// DATA
input [DATA_SIZE - 1:0] SIZE_W_IN;
input [DATA_SIZE - 1:0] V_IN;
output [DATA_SIZE - 1:0] V_OUT;

wire CLK;
wire RST;
wire START;
reg READY;
wire V_IN_ENABLE;
reg V_OUT_ENABLE;
wire [DATA_SIZE - 1:0] SIZE_W_IN;
wire [DATA_SIZE - 1:0] V_IN;
reg [DATA_SIZE - 1:0] V_OUT;


//---------------------------------------------------------------------
// Types
//---------------------------------------------------------------------
parameter [0:0]
  STARTER_STATE = 0,
  ENDER_STATE = 1;
  //---------------------------------------------------------------------
// Constants
//---------------------------------------------------------------------
parameter ZERO = ((0));
parameter ONE = ((1));  //---------------------------------------------------------------------
// Signals
//---------------------------------------------------------------------
// Finite State Machine
reg write_vector_ctrl_fsm_int;  // Internal Signals
reg [DATA_SIZE - 1:0] index_loop;

  //---------------------------------------------------------------------
  // Body
  //---------------------------------------------------------------------
  // v(t;k) = v^(t;k)
  always @(posedge CLK or posedge RST) begin
    if((RST == 1'b 0)) begin
      // Data Outputs
      V_OUT <= ZERO;
      // Control Outputs
      READY <= 1'b 0;
      // Assignations
      index_loop <= ZERO;
    end else begin
      case(write_vector_ctrl_fsm_int)
      STARTER_STATE : begin
        // STEP 0
        // Control Outputs
        READY <= 1'b 0;
        if((START == 1'b 1)) begin
          // Assignations
          index_loop <= ZERO;
          // FSM Control
          write_vector_ctrl_fsm_int <= ENDER_STATE;
        end
      end
      ENDER_STATE : begin
        // STEP 1
        if((V_IN_ENABLE == 1'b 1)) begin
          if((((index_loop)) == (((SIZE_W_IN)) - ((ONE))))) begin
            // Control Outputs
            READY <= 1'b 1;
            // FSM Control
            write_vector_ctrl_fsm_int <= STARTER_STATE;
          end
          else begin
            // Control Internal
            index_loop <= (((index_loop)) + ((ONE)));
          end
          // Data Outputs
          V_OUT <= V_IN;
          // Control Outputs
          V_OUT_ENABLE <= 1'b 1;
        end
        else begin
          // Control Outputs
          V_OUT_ENABLE <= 1'b 0;
        end
      end
      default : begin
        // FSM Control
        write_vector_ctrl_fsm_int <= STARTER_STATE;
      end
      endcase
    end
  end


endmodule
