--------------------------------------------------------------------------------
--                                            __ _      _     _               --
--                                           / _(_)    | |   | |              --
--                __ _ _   _  ___  ___ _ __ | |_ _  ___| | __| |              --
--               / _` | | | |/ _ \/ _ \ '_ \|  _| |/ _ \ |/ _` |              --
--              | (_| | |_| |  __/  __/ | | | | | |  __/ | (_| |              --
--               \__, |\__,_|\___|\___|_| |_|_| |_|\___|_|\__,_|              --
--                  | |                                                       --
--                  |_|                                                       --
--                                                                            --
--                                                                            --
--              Peripheral-NTM for MPSoC                                      --
--              Neural Turing Machine for MPSoC                               --
--                                                                            --
--------------------------------------------------------------------------------

-- Copyright (c) 2020-2021 by the author(s)
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
-- THE SOFTWARE.
--
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.ntm_math_pkg.all;

package dnc_core_pkg is

  -----------------------------------------------------------------------
  -- Constants
  -----------------------------------------------------------------------

  -----------------------------------------------------------------------
  -- Components
  -----------------------------------------------------------------------

  -----------------------------------------------------------------------
  -- MEMORY
  -----------------------------------------------------------------------

  component dnc_content_based_addressing is
    generic (
      I : integer := 64;
      J : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      K_IN_ENABLE : in std_logic; -- for j in 0 to J-1

      M_IN_I_ENABLE : in std_logic; -- for i in 0 to I-1
      M_IN_J_ENABLE : in std_logic; -- for j in 0 to J-1

      C_OUT_ENABLE : out std_logic; -- for i in 0 to I-1

      -- DATA
      K_IN    : in std_logic_vector(DATA_SIZE-1 downto 0);
      M_IN    : in std_logic_vector(DATA_SIZE-1 downto 0);
      BETA_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      C_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_allocation_weighting is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      PHI_IN_ENABLE : in std_logic; -- for j in 0 to N-1
      U_IN_ENABLE   : in std_logic; -- for j in 0 to N-1

      A_OUT_ENABLE : out std_logic; -- for j in 0 to N-1

      -- DATA
      PHI_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      U_IN   : in std_logic_vector(DATA_SIZE-1 downto 0);

      A_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_backward_weighting is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      L_IN_ENABLE : in std_logic; -- for j in 0 to N-1 (square matrix)

      W_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1 (read heads flow)
      W_IN_J_ENABLE : in std_logic; -- for j in 0 to N-1

      B_OUT_I_ENABLE : out std_logic; -- for i in 0 to R-1 (read heads flow)
      B_OUT_J_ENABLE : out std_logic; -- for j in 0 to N-1

      -- DATA
      L_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      W_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      B_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_forward_weighting is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      L_IN_ENABLE : in std_logic; -- for j in 0 to N-1 (square matrix)

      W_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1 (read heads flow)
      W_IN_J_ENABLE : in std_logic; -- for j in 0 to N-1

      F_OUT_I_ENABLE : out std_logic; -- for i in 0 to R-1 (read heads flow)
      F_OUT_J_ENABLE : out std_logic; -- for j in 0 to N-1

      -- DATA
      L_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      W_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      F_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_memory_matrix is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      M_IN_J_ENABLE : in std_logic; -- for j in 0 to N-1
      M_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1

      W_IN_J_ENABLE : in std_logic; -- for j in 0 to N-1
      V_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1
      E_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1

      M_OUT_J_ENABLE : out std_logic; -- for j in 0 to N-1
      M_OUT_K_ENABLE : out std_logic; -- for k in 0 to W-1

      -- DATA
      M_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      W_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      V_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      E_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      M_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_memory_retention_vector is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      F_IN_ENABLE : in std_logic; -- for i in 0 to R-1

      W_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1
      W_IN_J_ENABLE : in std_logic; -- for j in 0 to N-1

      PSI_OUT_ENABLE : out std_logic; -- for j in 0 to N-1

      -- DATA
      F_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      W_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      PSI_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_precedence_weighting is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      W_IN_ENABLE : in std_logic; -- for j in 0 to N-1
      P_IN_ENABLE : in std_logic; -- for j in 0 to N-1

      P_OUT_ENABLE : out std_logic; -- for j in 0 to N-1

      -- DATA
      W_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      P_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      P_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_read_content_weighting is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      K_IN_ENABLE : in std_logic; -- for k in 0 to W-1

      M_IN_J_ENABLE : in std_logic; -- for j in 0 to N-1
      M_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1

      C_OUT_ENABLE : out std_logic; -- for j in 0 to N-1

      -- DATA
      K_IN    : in std_logic_vector(DATA_SIZE-1 downto 0);
      M_IN    : in std_logic_vector(DATA_SIZE-1 downto 0);
      BETA_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      C_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_read_vectors is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      M_IN_J_ENABLE : in std_logic; -- for j in 0 to N-1
      M_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1

      W_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1 (read heads flow)
      W_IN_J_ENABLE : in std_logic; -- for j in 0 to N-1

      R_OUT_I_ENABLE : out std_logic; -- for i in 0 to R-1 (read heads flow)
      R_OUT_K_ENABLE : out std_logic; -- for k in 0 to W-1

        -- DATA
        M_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
        W_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      R_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_read_weighting is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      PI_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1
      PI_IN_P_ENABLE : in std_logic; -- for p in 0 to 2

      B_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1
      B_IN_J_ENABLE : in std_logic; -- for j in 0 to N-1

      C_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1
      C_IN_J_ENABLE : in std_logic; -- for j in 0 to N-1

      F_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1
      F_IN_J_ENABLE : in std_logic; -- for j in 0 to N-1

      W_OUT_I_ENABLE : out std_logic; -- for i in 0 to R-1
      W_OUT_J_ENABLE : out std_logic; -- for j in 0 to N-1

      -- DATA
      PI_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      B_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      C_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      F_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      W_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_sort_vector is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
     -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      U_IN_ENABLE : in std_logic; -- for j in 0 to N-1

      PHI_OUT_ENABLE : out std_logic; -- for j in 0 to N-1

      -- DATA
      U_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      PHI_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_temporal_link_matrix is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      L_IN_ENABLE : in std_logic; -- for j in 0 to N-1 (square matrix)
      W_IN_ENABLE : in std_logic; -- for j in 0 to N-1
      P_IN_ENABLE : in std_logic; -- for j in 0 to N-1

      L_OUT_ENABLE : out std_logic; -- for j in 0 to N-1

      -- DATA
      L_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      W_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      P_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      L_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_usage_vector is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      U_IN_ENABLE   : in std_logic; -- for j in 0 to N-1
      W_IN_ENABLE   : in std_logic; -- for j in 0 to N-1
      PSI_IN_ENABLE : in std_logic; -- for j in 0 to N-1

      U_OUT_ENABLE : out std_logic; -- for j in 0 to N-1

      -- DATA
      U_IN   : in std_logic_vector(DATA_SIZE-1 downto 0);
      W_IN   : in std_logic_vector(DATA_SIZE-1 downto 0);
      PSI_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      U_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_write_content_weighting is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      K_IN_ENABLE : in std_logic; -- for k in 0 to W-1

      M_IN_J_ENABLE : in std_logic; -- for j in 0 to N-1
      M_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1

      C_OUT_ENABLE : out std_logic; -- for j in 0 to N-1

      -- DATA
      K_IN    : in std_logic_vector(DATA_SIZE-1 downto 0);
      M_IN    : in std_logic_vector(DATA_SIZE-1 downto 0);
      BETA_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      C_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_write_weighting is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      A_IN_ENABLE : in std_logic; -- for j in 0 to N-1
      C_IN_ENABLE : in std_logic; -- for j in 0 to N-1

      W_OUT_ENABLE : out std_logic; -- for j in 0 to N-1

      -- DATA
      A_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      C_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      GA_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      GW_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      W_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_addressing is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      K_READ_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1
      K_READ_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1

      BETA_READ_IN_ENABLE : in std_logic; -- for i in 0 to R-1

      F_READ_IN_ENABLE : in std_logic; -- for i in 0 to R-1

      PI_READ_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1
      PI_READ_IN_P_ENABLE : in std_logic; -- for p in 0 to 2

      K_WRITE_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1
      E_WRITE_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1
      V_WRITE_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1

      -- DATA
      K_READ_IN    : in std_logic_vector(DATA_SIZE-1 downto 0);
      BETA_READ_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      F_READ_IN    : in std_logic_vector(DATA_SIZE-1 downto 0);
      PI_READ_IN   : in std_logic_vector(DATA_SIZE-1 downto 0);

      K_WRITE_IN    : in std_logic_vector(DATA_SIZE-1 downto 0);
      BETA_WRITE_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      E_WRITE_IN    : in std_logic_vector(DATA_SIZE-1 downto 0);
      V_WRITE_IN    : in std_logic_vector(DATA_SIZE-1 downto 0);
      GA_WRITE_IN   : in std_logic_vector(DATA_SIZE-1 downto 0);
      GW_WRITE_IN   : in std_logic_vector(DATA_SIZE-1 downto 0);

      R_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component dnc_addressing;

  -----------------------------------------------------------------------
  -- READ HEADS
  -----------------------------------------------------------------------

  component dnc_free_gates is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      F_IN_ENABLE : in std_logic; -- for i in 0 to R-1

      F_OUT_ENABLE : out std_logic; -- for i in 0 to R-1

      -- DATA
      F_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      F_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_read_keys is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      K_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1
      K_IN_J_ENABLE : in std_logic; -- for k in 0 to W-1

      K_OUT_I_ENABLE : out std_logic; -- for i in 0 to R-1
      K_OUT_J_ENABLE : out std_logic; -- for k in 0 to W-1

      -- DATA
      K_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      K_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_read_modes is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      PI_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1
      PI_IN_P_ENABLE : in std_logic; -- for p in 0 to 2

      PI_OUT_I_ENABLE : out std_logic; -- for i in 0 to R-1
      PI_OUT_P_ENABLE : out std_logic; -- for p in 0 to 2

      -- DATA
      PI_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      PI_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_read_strengths is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      BETA_IN_ENABLE : in std_logic; -- for i in 0 to R-1

      BETA_OUT_ENABLE : out std_logic; -- for i in 0 to R-1

      -- DATA
      BETA_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      BETA_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  -----------------------------------------------------------------------
  -- WRITE HEADS
  -----------------------------------------------------------------------

  component dnc_allocation_gate is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      -- DATA
      GA_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      GA_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_erase_vector is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      E_IN_ENABLE : in std_logic; -- for k in 0 to W-1

      E_OUT_ENABLE : out std_logic; -- for k in 0 to W-1

      -- DATA
      E_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      E_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_write_gate is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      -- DATA
      GW_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      GW_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_write_key is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      K_IN_ENABLE : in std_logic; -- for k in 0 to W-1

      K_OUT_ENABLE : out std_logic; -- for k in 0 to W-1

      -- DATA
      K_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      K_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_write_strength is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      -- DATA
      BETA_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      BETA_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_write_vector is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      V_IN_ENABLE : in std_logic; -- for k in 0 to W-1

      V_OUT_ENABLE : out std_logic; -- for k in 0 to W-1

      -- DATA
      V_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      V_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  -----------------------------------------------------------------------
  -- TOP
  -----------------------------------------------------------------------

  component dnc_top is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      X_IN_ENABLE : in std_logic; -- for x in 0 to X-1

      Y_OUT_ENABLE : out std_logic; -- for y in 0 to Y-1

      -- DATA
      X_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      Y_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_output_vector is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      K_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1
      K_IN_Y_ENABLE : in std_logic; -- for y in 0 to Y-1
      K_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1

      R_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1
      R_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1

      NU_IN_ENABLE : in std_logic; -- for y in 0 to Y-1

      Y_OUT_ENABLE : in std_logic; -- for y in 0 to Y-1

      -- DATA
      K_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      R_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      NU_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      Y_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_controller_output_vector is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      U_IN_Y_ENABLE : in std_logic; -- for y in 0 to Y-1
      U_IN_L_ENABLE : in std_logic; -- for l in 0 to L-1

      H_IN_ENABLE : in std_logic; -- for l in 0 to L-1

      NU_ENABLE_OUT : out std_logic; -- for j in 0 to Y-1

      -- DATA
      U_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      H_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      NU_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_read_interface_vector is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      -- Read Key
      WK_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1
      WK_IN_L_ENABLE : in std_logic; -- for l in 0 to L-1
      WK_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1

      K_OUT_I_ENABLE : in std_logic; -- for i in 0 to R-1
      K_OUT_K_ENABLE : in std_logic; -- for k in 0 to W-1

      -- Read Strength
      WBETA_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1
      WBETA_IN_L_ENABLE : in std_logic; -- for l in 0 to L-1

      BETA_OUT_ENABLE : in std_logic; -- for i in 0 to R-1

      -- Free Gate
      WF_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1
      WF_IN_L_ENABLE : in std_logic; -- for l in 0 to L-1

      F_OUT_ENABLE : in std_logic; -- for i in 0 to R-1

      -- Read Mode
      WPI_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1
      WPI_IN_L_ENABLE : in std_logic; -- for l in 0 to L-1
      WPI_IN_P_ENABLE : in std_logic; -- for p in 0 to 2

      PI_OUT_I_ENABLE : in std_logic; -- for i in 0 to R-1
      PI_OUT_P_ENABLE : in std_logic; -- for p in 0 to 2

      -- Hidden State
      H_IN_ENABLE : in std_logiC; -- for l in 0 to L-1

      -- DATA
      WK_IN    : in std_logic_vector(DATA_SIZE-1 downto 0);
      WBETA_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      WF_IN    : in std_logic_vector(DATA_SIZE-1 downto 0);
      WPI_IN   : in std_logic_vector(DATA_SIZE-1 downto 0);

      H_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      K_OUT    : out std_logic_vector(DATA_SIZE-1 downto 0);
      BETA_OUT : out std_logic_vector(DATA_SIZE-1 downto 0);
      F_OUT    : out std_logic_vector(DATA_SIZE-1 downto 0);
      PI_OUT   : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component dnc_write_interface_vector is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;
      R : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      -- Write Key
      WK_IN_L_ENABLE : in std_logic; -- for l in 0 to L-1
      WK_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1

      K_OUT_ENABLE : out std_logic; -- for k in 0 to W-1

      -- Write Strength
      WBETA_IN_ENABLE : in std_logic; -- for l in 0 to L-1

      -- Erase Vector
      WE_IN_L_ENABLE : in std_logic; -- for l in 0 to L-1
      WE_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1

      E_OUT_ENABLE : out std_logic; -- for k in 0 to W-1

      -- Write Vector
      WV_IN_L_ENABLE : in std_logic; -- for l in 0 to L-1
      WV_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1

      V_OUT_ENABLE : out std_logic; -- for k in 0 to W-1

      -- Allocation Gate
      WGA_IN_ENABLE : in std_logic; -- for l in 0 to L-1

      -- Write Gate
      WGW_IN_ENABLE : in std_logic; -- for l in 0 to L-1

      -- Hidden State
      H_IN_ENABLE : in std_logic; -- for l in 0 to L-1

      -- DATA
      WK_IN    : in std_logic_vector(DATA_SIZE-1 downto 0);
      WBETA_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      WE_IN    : in std_logic_vector(DATA_SIZE-1 downto 0);
      WV_IN    : in std_logic_vector(DATA_SIZE-1 downto 0);
      WGA_IN   : in std_logic_vector(DATA_SIZE-1 downto 0);
      WGW_IN   : in std_logic_vector(DATA_SIZE-1 downto 0);

      H_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      K_OUT    : out std_logic_vector(DATA_SIZE-1 downto 0);
      BETA_OUT : out std_logic_vector(DATA_SIZE-1 downto 0);
      E_OUT    : out std_logic_vector(DATA_SIZE-1 downto 0);
      V_OUT    : out std_logic_vector(DATA_SIZE-1 downto 0);
      GA_OUT   : out std_logic_vector(DATA_SIZE-1 downto 0);
      GW_OUT   : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

end dnc_core_pkg;
