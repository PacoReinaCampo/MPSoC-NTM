////////////////////////////////////////////////////////////////////////////////
//                                            __ _      _     _               //
//                                           / _(_)    | |   | |              //
//                __ _ _   _  ___  ___ _ __ | |_ _  ___| | __| |              //
//               / _` | | | |/ _ \/ _ \ '_ \|  _| |/ _ \ |/ _` |              //
//              | (_| | |_| |  __/  __/ | | | | | |  __/ | (_| |              //
//               \__, |\__,_|\___|\___|_| |_|_| |_|\___|_|\__,_|              //
//                  | |                                                       //
//                  |_|                                                       //
//                                                                            //
//                                                                            //
//              Peripheral-NTM for MPSoC                                      //
//              Neural Turing Machine for MPSoC                               //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2020-2021 by the author(s)
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
////////////////////////////////////////////////////////////////////////////////
// Author(s):
//   Paco Reina Campo <pacoreinacampo@queenfield.tech>

package ntm_function_pkg;

  ///////////////////////////////////////////////////////////////////////
  // Types
  ///////////////////////////////////////////////////////////////////////

  ///////////////////////////////////////////////////////////////////////
  // Constants
  ///////////////////////////////////////////////////////////////////////

  // SYSTEM-SIZE
  parameter DATA_SIZE=128;
  parameter CONTROL_SIZE=64;

  parameter X=64;
  parameter Y=64;
  parameter N=64;
  parameter W=64;
  parameter L=64;
  parameter R=64;

  // SCALAR-FUNCTIONALITY
  parameter STIMULUS_NTM_SCALAR_CONVOLUTION_TEST=0;
  parameter STIMULUS_NTM_SCALAR_COSINE_SIMILARITY_TEST=0;
  parameter STIMULUS_NTM_SCALAR_COSH_TEST=0;
  parameter STIMULUS_NTM_SCALAR_SINH_TEST=0;
  parameter STIMULUS_NTM_SCALAR_TANH_TEST=0;
  parameter STIMULUS_NTM_SCALAR_LOGISTIC_TEST=0;
  parameter STIMULUS_NTM_SCALAR_SOFTMAX_TEST=0;
  parameter STIMULUS_NTM_SCALAR_ONE_CONTROLPLUS_TEST=0;
  parameter STIMULUS_NTM_SCALAR_SUMMATION_TEST=0;
  parameter STIMULUS_NTM_SCALAR_CONVOLUTION_CASE_0=0;
  parameter STIMULUS_NTM_SCALAR_COSINE_SIMILARITY_CASE_0=0;
  parameter STIMULUS_NTM_SCALAR_COSH_CASE_0=0;
  parameter STIMULUS_NTM_SCALAR_SINH_CASE_0=0;
  parameter STIMULUS_NTM_SCALAR_TANH_CASE_0=0;
  parameter STIMULUS_NTM_SCALAR_LOGISTIC_CASE_0=0;
  parameter STIMULUS_NTM_SCALAR_SOFTMAX_CASE_0=0;
  parameter STIMULUS_NTM_SCALAR_ONE_CONTROLPLUS_CASE_0=0;
  parameter STIMULUS_NTM_SCALAR_SUMMATION_CASE_0=0;
  parameter STIMULUS_NTM_SCALAR_CONVOLUTION_CASE_1=0;
  parameter STIMULUS_NTM_SCALAR_COSINE_SIMILARITY_CASE_1=0;
  parameter STIMULUS_NTM_SCALAR_COSH_CASE_1=0;
  parameter STIMULUS_NTM_SCALAR_SINH_CASE_1=0;
  parameter STIMULUS_NTM_SCALAR_TANH_CASE_1=0;
  parameter STIMULUS_NTM_SCALAR_LOGISTIC_CASE_1=0;
  parameter STIMULUS_NTM_SCALAR_SOFTMAX_CASE_1=0;
  parameter STIMULUS_NTM_SCALAR_ONE_CONTROLPLUS_CASE_1=0;
  parameter STIMULUS_NTM_SCALAR_SUMMATION_CASE_1=0;

  // VECTOR-FUNCTIONALITY
  parameter STIMULUS_NTM_VECTOR_CONVOLUTION_TEST=0;
  parameter STIMULUS_NTM_VECTOR_COSINE_SIMILARITY_TEST=0;
  parameter STIMULUS_NTM_VECTOR_COSH_TEST=0;
  parameter STIMULUS_NTM_VECTOR_SINH_TEST=0;
  parameter STIMULUS_NTM_VECTOR_TANH_TEST=0;
  parameter STIMULUS_NTM_VECTOR_LOGISTIC_TEST=0;
  parameter STIMULUS_NTM_VECTOR_SOFTMAX_TEST=0;
  parameter STIMULUS_NTM_VECTOR_ONE_CONTROLPLUS_TEST=0;
  parameter STIMULUS_NTM_VECTOR_SUMMATION_TEST=0;
  parameter STIMULUS_NTM_VECTOR_CONVOLUTION_CASE_0=0;
  parameter STIMULUS_NTM_VECTOR_COSINE_SIMILARITY_CASE_0=0;
  parameter STIMULUS_NTM_VECTOR_COSH_CASE_0=0;
  parameter STIMULUS_NTM_VECTOR_SINH_CASE_0=0;
  parameter STIMULUS_NTM_VECTOR_TANH_CASE_0=0;
  parameter STIMULUS_NTM_VECTOR_LOGISTIC_CASE_0=0;
  parameter STIMULUS_NTM_VECTOR_SOFTMAX_CASE_0=0;
  parameter STIMULUS_NTM_VECTOR_ONE_CONTROLPLUS_CASE_0=0;
  parameter STIMULUS_NTM_VECTOR_SUMMATION_CASE_0=0;
  parameter STIMULUS_NTM_VECTOR_CONVOLUTION_CASE_1=0;
  parameter STIMULUS_NTM_VECTOR_COSINE_SIMILARITY_CASE_1=0;
  parameter STIMULUS_NTM_VECTOR_COSH_CASE_1=0;
  parameter STIMULUS_NTM_VECTOR_SINH_CASE_1=0;
  parameter STIMULUS_NTM_VECTOR_TANH_CASE_1=0;
  parameter STIMULUS_NTM_VECTOR_LOGISTIC_CASE_1=0;
  parameter STIMULUS_NTM_VECTOR_SOFTMAX_CASE_1=0;
  parameter STIMULUS_NTM_VECTOR_ONE_CONTROLPLUS_CASE_1=0;
  parameter STIMULUS_NTM_VECTOR_SUMMATION_CASE_1=0;

  // MATRIX-FUNCTIONALITY
  parameter STIMULUS_NTM_MATRIX_CONVOLUTION_TEST=0;
  parameter STIMULUS_NTM_MATRIX_COSINE_SIMILARITY_TEST=0;
  parameter STIMULUS_NTM_MATRIX_COSH_TEST=0;
  parameter STIMULUS_NTM_MATRIX_SINH_TEST=0;
  parameter STIMULUS_NTM_MATRIX_TANH_TEST=0;
  parameter STIMULUS_NTM_MATRIX_LOGISTIC_TEST=0;
  parameter STIMULUS_NTM_MATRIX_SOFTMAX_TEST=0;
  parameter STIMULUS_NTM_MATRIX_ONE_CONTROLPLUS_TEST=0;
  parameter STIMULUS_NTM_MATRIX_SUMMATION_TEST=0;
  parameter STIMULUS_NTM_MATRIX_CONVOLUTION_CASE_0=0;
  parameter STIMULUS_NTM_MATRIX_COSINE_SIMILARITY_CASE_0=0;
  parameter STIMULUS_NTM_MATRIX_COSH_CASE_0=0;
  parameter STIMULUS_NTM_MATRIX_SINH_CASE_0=0;
  parameter STIMULUS_NTM_MATRIX_TANH_CASE_0=0;
  parameter STIMULUS_NTM_MATRIX_LOGISTIC_CASE_0=0;
  parameter STIMULUS_NTM_MATRIX_SOFTMAX_CASE_0=0;
  parameter STIMULUS_NTM_MATRIX_ONE_CONTROLPLUS_CASE_0=0;
  parameter STIMULUS_NTM_MATRIX_SUMMATION_CASE_0=0;
  parameter STIMULUS_NTM_MATRIX_CONVOLUTION_CASE_1=0;
  parameter STIMULUS_NTM_MATRIX_COSINE_SIMILARITY_CASE_1=0;
  parameter STIMULUS_NTM_MATRIX_COSH_CASE_1=0;
  parameter STIMULUS_NTM_MATRIX_SINH_CASE_1=0;
  parameter STIMULUS_NTM_MATRIX_TANH_CASE_1=0;
  parameter STIMULUS_NTM_MATRIX_LOGISTIC_CASE_1=0;
  parameter STIMULUS_NTM_MATRIX_SOFTMAX_CASE_1=0;
  parameter STIMULUS_NTM_MATRIX_ONE_CONTROLPLUS_CASE_1=0;
  parameter STIMULUS_NTM_MATRIX_SUMMATION_CASE_1=0;

  ///////////////////////////////////////////////////////////////////////
  // Signals
  ///////////////////////////////////////////////////////////////////////

endpackage
