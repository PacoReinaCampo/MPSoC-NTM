--------------------------------------------------------------------------------
--                                            __ _      _     _               --
--                                           / _(_)    | |   | |              --
--                __ _ _   _  ___  ___ _ __ | |_ _  ___| | __| |              --
--               / _` | | | |/ _ \/ _ \ '_ \|  _| |/ _ \ |/ _` |              --
--              | (_| | |_| |  __/  __/ | | | | | |  __/ | (_| |              --
--               \__, |\__,_|\___|\___|_| |_|_| |_|\___|_|\__,_|              --
--                  | |                                                       --
--                  |_|                                                       --
--                                                                            --
--                                                                            --
--              Peripheral-NTM for MPSoC                                      --
--              Neural Turing Machine for MPSoC                               --
--                                                                            --
--------------------------------------------------------------------------------

-- Copyright (c) 2020-2021 by the author(s)
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
-- THE SOFTWARE.
--
--------------------------------------------------------------------------------
-- Author(s):
--   Paco Reina Campo <pacoreinacampo@queenfield.tech>

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.ntm_math_pkg.all;

entity ntm_scalar_adder is
  generic (
    DATA_SIZE    : integer := 128;
    CONTROL_SIZE : integer := 64
    );
  port (
    -- GLOBAL
    CLK : in std_logic;
    RST : in std_logic;

    -- CONTROL
    START : in  std_logic;
    READY : out std_logic;

    OPERATION : in std_logic;

    -- DATA
    DATA_A_IN : in  std_logic_vector(DATA_SIZE-1 downto 0);
    DATA_B_IN : in  std_logic_vector(DATA_SIZE-1 downto 0);

    DATA_OUT     : out std_logic_vector(DATA_SIZE-1 downto 0);
    OVERFLOW_OUT : out std_logic
    );
end entity;

architecture ntm_scalar_adder_architecture of ntm_scalar_adder is

  -----------------------------------------------------------------------
  -- Types
  -----------------------------------------------------------------------

  type adder_ctrl_fsm is (
    STARTER_STATE,                      -- STEP 0
    ARITHMETIC_STATE,                   -- STEP 1
    ADAPTATION_STATE,                   -- STEP 2
    NORMALIZATION_STATE,                -- STEP 3
    ENDER_STATE                         -- STEP 4
    );

  -----------------------------------------------------------------------
  -- Constants
  -----------------------------------------------------------------------

  constant EXPONENT_SIZE : integer := 15;
  constant MANTISSA_SIZE : integer := 112;

  constant ZERO_EXPONENT  : std_logic_vector(EXPONENT_SIZE-1 downto 0) := std_logic_vector(to_unsigned(0, EXPONENT_SIZE));
  constant ONE_EXPONENT   : std_logic_vector(EXPONENT_SIZE-1 downto 0) := std_logic_vector(to_unsigned(1, EXPONENT_SIZE));
  constant TWO_EXPONENT   : std_logic_vector(EXPONENT_SIZE-1 downto 0) := std_logic_vector(to_unsigned(2, EXPONENT_SIZE));
  constant THREE_EXPONENT : std_logic_vector(EXPONENT_SIZE-1 downto 0) := std_logic_vector(to_unsigned(3, EXPONENT_SIZE));

  constant ZERO_MANTISSA  : std_logic_vector(MANTISSA_SIZE-1 downto 0) := std_logic_vector(to_unsigned(0, MANTISSA_SIZE));
  constant ONE_MANTISSA   : std_logic_vector(MANTISSA_SIZE-1 downto 0) := std_logic_vector(to_unsigned(1, MANTISSA_SIZE));
  constant TWO_MANTISSA   : std_logic_vector(MANTISSA_SIZE-1 downto 0) := std_logic_vector(to_unsigned(2, MANTISSA_SIZE));
  constant THREE_MANTISSA : std_logic_vector(MANTISSA_SIZE-1 downto 0) := std_logic_vector(to_unsigned(3, MANTISSA_SIZE));

  constant ZERO_CONTROL  : std_logic_vector(CONTROL_SIZE-1 downto 0) := std_logic_vector(to_unsigned(0, CONTROL_SIZE));
  constant ONE_CONTROL   : std_logic_vector(CONTROL_SIZE-1 downto 0) := std_logic_vector(to_unsigned(1, CONTROL_SIZE));
  constant TWO_CONTROL   : std_logic_vector(CONTROL_SIZE-1 downto 0) := std_logic_vector(to_unsigned(2, CONTROL_SIZE));
  constant THREE_CONTROL : std_logic_vector(CONTROL_SIZE-1 downto 0) := std_logic_vector(to_unsigned(3, CONTROL_SIZE));

  constant ZERO_DATA  : std_logic_vector(DATA_SIZE-1 downto 0) := std_logic_vector(to_unsigned(0, DATA_SIZE));
  constant ONE_DATA   : std_logic_vector(DATA_SIZE-1 downto 0) := std_logic_vector(to_unsigned(1, DATA_SIZE));
  constant TWO_DATA   : std_logic_vector(DATA_SIZE-1 downto 0) := std_logic_vector(to_unsigned(2, DATA_SIZE));
  constant THREE_DATA : std_logic_vector(DATA_SIZE-1 downto 0) := std_logic_vector(to_unsigned(3, DATA_SIZE));

  constant FULL  : std_logic_vector(DATA_SIZE-1 downto 0) := (others => '1');
  constant EMPTY : std_logic_vector(DATA_SIZE-1 downto 0) := (others => '0');

  constant FULL_EXPONENT  : std_logic_vector(EXPONENT_SIZE-1 downto 0) := (others => '1');
  constant EMPTY_EXPONENT : std_logic_vector(EXPONENT_SIZE-1 downto 0) := (others => '0');

  constant FULL_MANTISSA  : std_logic_vector(MANTISSA_SIZE-1 downto 0) := (others => '1');
  constant EMPTY_MANTISSA : std_logic_vector(MANTISSA_SIZE-1 downto 0) := (others => '0');

  constant EULER : std_logic_vector(DATA_SIZE-1 downto 0) := (others => '0');

  constant BIAS : std_logic_vector(EXPONENT_SIZE-1 downto 0) := std_logic_vector(to_unsigned(2**(EXPONENT_SIZE-1)-1, EXPONENT_SIZE));

  -----------------------------------------------------------------------
  -- Signals
  -----------------------------------------------------------------------

  -- Finite State Machine
  signal adder_ctrl_fsm_int : adder_ctrl_fsm;

  -- EXPONENT SCALAR ADDER
  -- CONTROL
  signal start_exponent_scalar_adder : std_logic;
  signal ready_exponent_scalar_adder : std_logic;

  signal operation_exponent_scalar_adder : std_logic;

  -- DATA
  signal data_a_in_exponent_scalar_adder : std_logic_vector(EXPONENT_SIZE-1 downto 0);
  signal data_b_in_exponent_scalar_adder : std_logic_vector(EXPONENT_SIZE-1 downto 0);

  signal data_out_exponent_scalar_adder     : std_logic_vector(EXPONENT_SIZE-1 downto 0);
  signal overflow_out_exponent_scalar_adder : std_logic;

  -- MANTISSA SCALAR ADDER
  -- CONTROL
  signal start_mantissa_scalar_adder : std_logic;
  signal ready_mantissa_scalar_adder : std_logic;

  signal operation_mantissa_scalar_adder : std_logic;

  -- DATA
  signal data_a_in_mantissa_scalar_adder : std_logic_vector(MANTISSA_SIZE-1 downto 0);
  signal data_b_in_mantissa_scalar_adder : std_logic_vector(MANTISSA_SIZE-1 downto 0);

  signal data_out_mantissa_scalar_adder     : std_logic_vector(MANTISSA_SIZE-1 downto 0);
  signal overflow_out_mantissa_scalar_adder : std_logic;

  -- OUTPUT
  signal sign_int_scalar_adder : std_logic;

  signal exponent_int_scalar_adder : std_logic_vector(EXPONENT_SIZE-1 downto 0);
  signal mantissa_int_scalar_adder : std_logic_vector(MANTISSA_SIZE-1 downto 0);

begin

  -----------------------------------------------------------------------
  -- Body
  -----------------------------------------------------------------------

  -- DATA_OUT = DATA_A_IN ± DATA_B_IN = M_A_IN · 2^(E_A_IN) ± M_B_IN · 2^(E_B_IN)

  -- CONTROL
  ctrl_fsm : process(CLK, RST)
  begin
    if (RST = '0') then
      -- Data Outputs
      DATA_OUT <= ZERO_DATA;

      -- Control Outputs
      READY <= '0';

      -- Control Internal
      start_exponent_scalar_adder <= '0';
      start_mantissa_scalar_adder <= '0';

      operation_exponent_scalar_adder <= '0';
      operation_mantissa_scalar_adder <= '0';

      -- Data Internal
      data_a_in_exponent_scalar_adder <= ZERO_EXPONENT;
      data_b_in_exponent_scalar_adder <= ZERO_EXPONENT;

      data_a_in_mantissa_scalar_adder <= ZERO_MANTISSA;
      data_b_in_mantissa_scalar_adder <= ZERO_MANTISSA;

      sign_int_scalar_adder <= '0';

      exponent_int_scalar_adder <= ZERO_EXPONENT;
      mantissa_int_scalar_adder <= ZERO_MANTISSA;

    elsif (rising_edge(CLK)) then

      case adder_ctrl_fsm_int is
        when STARTER_STATE =>  -- STEP 0
          -- Control Outputs
          READY <= '0';

          if (START = '1') then
            -- Control Internal
            start_exponent_scalar_adder <= '1';
            start_mantissa_scalar_adder <= '1';

            operation_exponent_scalar_adder <= '0';
            operation_mantissa_scalar_adder <= '0';

            -- Data Internal
            sign_int_scalar_adder <= DATA_A_IN(DATA_SIZE-1) xor DATA_B_IN(DATA_SIZE-1);

            data_a_in_exponent_scalar_adder <= DATA_A_IN(DATA_SIZE-2 downto MANTISSA_SIZE);
            data_b_in_exponent_scalar_adder <= DATA_B_IN(DATA_SIZE-2 downto MANTISSA_SIZE);

            data_a_in_mantissa_scalar_adder <= DATA_A_IN(MANTISSA_SIZE-1 downto 0);
            data_b_in_mantissa_scalar_adder <= DATA_B_IN(MANTISSA_SIZE-1 downto 0);

            -- FSM Control
            adder_ctrl_fsm_int <= ARITHMETIC_STATE;
          end if;

        when ARITHMETIC_STATE =>  -- STEP 1

          if (ready_exponent_scalar_adder = '1') then
            -- Data Outputs
            exponent_int_scalar_adder <= data_out_exponent_scalar_adder;
          else
            -- Control Internal
            start_exponent_scalar_adder <= '0';
          end if;

          if (ready_mantissa_scalar_adder = '1') then
            -- Data Outputs
            mantissa_int_scalar_adder <= data_out_mantissa_scalar_adder;
          else
            -- Control Internal
            start_mantissa_scalar_adder <= '0';
          end if;

        when ADAPTATION_STATE =>  -- STEP 2

          if (exponent_int_scalar_adder(EXPONENT_SIZE-1) = '1') then
            -- Data Outputs
            exponent_int_scalar_adder <= std_logic_vector(unsigned(exponent_int_scalar_adder) - unsigned(ONE_EXPONENT));
            mantissa_int_scalar_adder <= std_logic_vector(unsigned(mantissa_int_scalar_adder) sll 1);
          end if;

        when NORMALIZATION_STATE =>  -- STEP 3

        when ENDER_STATE =>  -- STEP 4

          -- Control Outputs
          READY <= '1';

          -- Data Outputs
          DATA_OUT <= sign_int_scalar_adder & exponent_int_scalar_adder & mantissa_int_scalar_adder;

        when others =>
          -- FSM Control
          adder_ctrl_fsm_int <= STARTER_STATE;
      end case;
    end if;
  end process;

  -- EXPONENT SCALAR ADDER
  exponent_scalar_adder : ntm_scalar_integer_adder
    generic map (
      DATA_SIZE    => EXPONENT_SIZE,
      CONTROL_SIZE => CONTROL_SIZE
      )
    port map (
      -- GLOBAL
      CLK => CLK,
      RST => RST,

      -- CONTROL
      START => start_exponent_scalar_adder,
      READY => ready_exponent_scalar_adder,

      OPERATION => operation_exponent_scalar_adder,

      -- DATA
      DATA_A_IN => data_a_in_exponent_scalar_adder,
      DATA_B_IN => data_b_in_exponent_scalar_adder,

      DATA_OUT     => data_out_exponent_scalar_adder,
      OVERFLOW_OUT => overflow_out_exponent_scalar_adder
      );

  -- MANTISSA SCALAR ADDER
  mantissa_scalar_adder : ntm_scalar_integer_adder
    generic map (
      DATA_SIZE    => MANTISSA_SIZE,
      CONTROL_SIZE => CONTROL_SIZE
      )
    port map (
      -- GLOBAL
      CLK => CLK,
      RST => RST,

      -- CONTROL
      START => start_mantissa_scalar_adder,
      READY => ready_mantissa_scalar_adder,

      OPERATION => operation_mantissa_scalar_adder,

      -- DATA
      DATA_A_IN => data_a_in_mantissa_scalar_adder,
      DATA_B_IN => data_b_in_mantissa_scalar_adder,

      DATA_OUT     => data_out_mantissa_scalar_adder,
      OVERFLOW_OUT => overflow_out_mantissa_scalar_adder
      );

end architecture;
