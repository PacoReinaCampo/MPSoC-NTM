--------------------------------------------------------------------------------
--                                            __ _      _     _               --
--                                           / _(_)    | |   | |              --
--                __ _ _   _  ___  ___ _ __ | |_ _  ___| | __| |              --
--               / _` | | | |/ _ \/ _ \ '_ \|  _| |/ _ \ |/ _` |              --
--              | (_| | |_| |  __/  __/ | | | | | |  __/ | (_| |              --
--               \__, |\__,_|\___|\___|_| |_|_| |_|\___|_|\__,_|              --
--                  | |                                                       --
--                  |_|                                                       --
--                                                                            --
--                                                                            --
--              Peripheral-NTM for MPSoC                                      --
--              Neural Turing Machine for MPSoC                               --
--                                                                            --
--------------------------------------------------------------------------------

-- Copyright (c) 2020-2021 by the author(s)
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
-- THE SOFTWARE.
--
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.ntm_math_pkg.all;
use work.ntm_function_pkg.all;

entity ntm_function_testbench is
  generic (
    -- SYSTEM-SIZE
    DATA_SIZE    : integer := 128;
    CONTROL_SIZE : integer := 64;

    X : std_logic_vector(DATA_SIZE-1 downto 0) := std_logic_vector(to_unsigned(64, DATA_SIZE));  -- x in 0 to X-1
    Y : std_logic_vector(DATA_SIZE-1 downto 0) := std_logic_vector(to_unsigned(64, DATA_SIZE));  -- y in 0 to Y-1
    N : std_logic_vector(DATA_SIZE-1 downto 0) := std_logic_vector(to_unsigned(64, DATA_SIZE));  -- j in 0 to N-1
    W : std_logic_vector(DATA_SIZE-1 downto 0) := std_logic_vector(to_unsigned(64, DATA_SIZE));  -- k in 0 to W-1
    L : std_logic_vector(DATA_SIZE-1 downto 0) := std_logic_vector(to_unsigned(64, DATA_SIZE));  -- l in 0 to L-1
    R : std_logic_vector(DATA_SIZE-1 downto 0) := std_logic_vector(to_unsigned(64, DATA_SIZE));  -- i in 0 to R-1

    -- SCALAR-FUNCTIONALITY
    ENABLE_NTM_SCALAR_COSH_TEST          : boolean := false;
    ENABLE_NTM_SCALAR_EXPONENTIATOR_TEST : boolean := false;
    ENABLE_NTM_SCALAR_LOGARITHM_TEST     : boolean := false;
    ENABLE_NTM_SCALAR_LOGISTIC_TEST      : boolean := false;
    ENABLE_NTM_SCALAR_ONEPLUS_TEST       : boolean := false;
    ENABLE_NTM_SCALAR_SINH_TEST          : boolean := false;
    ENABLE_NTM_SCALAR_TANH_TEST          : boolean := false;

    ENABLE_NTM_SCALAR_COSH_CASE_0          : boolean := false;
    ENABLE_NTM_SCALAR_EXPONENTIATOR_CASE_0 : boolean := false;
    ENABLE_NTM_SCALAR_LOGARITHM_CASE_0     : boolean := false;
    ENABLE_NTM_SCALAR_LOGISTIC_CASE_0      : boolean := false;
    ENABLE_NTM_SCALAR_ONEPLUS_CASE_0       : boolean := false;
    ENABLE_NTM_SCALAR_SINH_CASE_0          : boolean := false;
    ENABLE_NTM_SCALAR_TANH_CASE_0          : boolean := false;

    ENABLE_NTM_SCALAR_COSH_CASE_1          : boolean := false;
    ENABLE_NTM_SCALAR_EXPONENTIATOR_CASE_1 : boolean := false;
    ENABLE_NTM_SCALAR_LOGARITHM_CASE_1     : boolean := false;
    ENABLE_NTM_SCALAR_LOGISTIC_CASE_1      : boolean := false;
    ENABLE_NTM_SCALAR_ONEPLUS_CASE_1       : boolean := false;
    ENABLE_NTM_SCALAR_SINH_CASE_1          : boolean := false;
    ENABLE_NTM_SCALAR_TANH_CASE_1          : boolean := false;

    -- VECTOR-FUNCTIONALITY
    ENABLE_NTM_VECTOR_COSH_TEST          : boolean := false;
    ENABLE_NTM_VECTOR_EXPONENTIATOR_TEST : boolean := false;
    ENABLE_NTM_VECTOR_LOGARITHM_TEST     : boolean := false;
    ENABLE_NTM_VECTOR_LOGISTIC_TEST      : boolean := false;
    ENABLE_NTM_VECTOR_ONEPLUS_TEST       : boolean := false;
    ENABLE_NTM_VECTOR_SINH_TEST          : boolean := false;
    ENABLE_NTM_VECTOR_TANH_TEST          : boolean := false;

    ENABLE_NTM_VECTOR_COSH_CASE_0          : boolean := false;
    ENABLE_NTM_VECTOR_EXPONENTIATOR_CASE_0 : boolean := false;
    ENABLE_NTM_VECTOR_LOGARITHM_CASE_0     : boolean := false;
    ENABLE_NTM_VECTOR_LOGISTIC_CASE_0      : boolean := false;
    ENABLE_NTM_VECTOR_ONEPLUS_CASE_0       : boolean := false;
    ENABLE_NTM_VECTOR_SINH_CASE_0          : boolean := false;
    ENABLE_NTM_VECTOR_TANH_CASE_0          : boolean := false;

    ENABLE_NTM_VECTOR_COSH_CASE_1          : boolean := false;
    ENABLE_NTM_VECTOR_EXPONENTIATOR_CASE_1 : boolean := false;
    ENABLE_NTM_VECTOR_LOGARITHM_CASE_1     : boolean := false;
    ENABLE_NTM_VECTOR_LOGISTIC_CASE_1      : boolean := false;
    ENABLE_NTM_VECTOR_ONEPLUS_CASE_1       : boolean := false;
    ENABLE_NTM_VECTOR_SINH_CASE_1          : boolean := false;
    ENABLE_NTM_VECTOR_TANH_CASE_1          : boolean := false;

    -- MATRIX-FUNCTIONALITY
    ENABLE_NTM_MATRIX_COSH_TEST          : boolean := false;
    ENABLE_NTM_MATRIX_EXPONENTIATOR_TEST : boolean := false;
    ENABLE_NTM_MATRIX_LOGARITHM_TEST     : boolean := false;
    ENABLE_NTM_MATRIX_LOGISTIC_TEST      : boolean := false;
    ENABLE_NTM_MATRIX_ONEPLUS_TEST       : boolean := false;
    ENABLE_NTM_MATRIX_SINH_TEST          : boolean := false;
    ENABLE_NTM_MATRIX_TANH_TEST          : boolean := false;

    ENABLE_NTM_MATRIX_COSH_CASE_0          : boolean := false;
    ENABLE_NTM_MATRIX_EXPONENTIATOR_CASE_0 : boolean := false;
    ENABLE_NTM_MATRIX_LOGARITHM_CASE_0     : boolean := false;
    ENABLE_NTM_MATRIX_LOGISTIC_CASE_0      : boolean := false;
    ENABLE_NTM_MATRIX_ONEPLUS_CASE_0       : boolean := false;
    ENABLE_NTM_MATRIX_SINH_CASE_0          : boolean := false;
    ENABLE_NTM_MATRIX_TANH_CASE_0          : boolean := false;

    ENABLE_NTM_MATRIX_COSH_CASE_1          : boolean := false;
    ENABLE_NTM_MATRIX_EXPONENTIATOR_CASE_1 : boolean := false;
    ENABLE_NTM_MATRIX_LOGARITHM_CASE_1     : boolean := false;
    ENABLE_NTM_MATRIX_LOGISTIC_CASE_1      : boolean := false;
    ENABLE_NTM_MATRIX_ONEPLUS_CASE_1       : boolean := false;
    ENABLE_NTM_MATRIX_SINH_CASE_1          : boolean := false;
    ENABLE_NTM_MATRIX_TANH_CASE_1          : boolean := false
    );
end ntm_function_testbench;

architecture ntm_function_testbench_architecture of ntm_function_testbench is

  -----------------------------------------------------------------------
  -- Signals
  -----------------------------------------------------------------------

  -- GLOBAL
  signal CLK : std_logic;
  signal RST : std_logic;

  -----------------------------------------------------------------------
  -- SCALAR
  -----------------------------------------------------------------------

  -- SCALAR COSH
  -- CONTROL
  signal start_scalar_cosh : std_logic;
  signal ready_scalar_cosh : std_logic;

  -- DATA
  signal data_in_scalar_cosh  : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_scalar_cosh : std_logic_vector(DATA_SIZE-1 downto 0);

  -- CONTROL
  signal start_scalar_cosine_similarity : std_logic;
  signal ready_scalar_cosine_similarity : std_logic;

  signal data_a_in_enable_scalar_cosine_similarity : std_logic;
  signal data_b_in_enable_scalar_cosine_similarity : std_logic;

  signal data_out_enable_scalar_cosine_similarity : std_logic;

  -- DATA
  signal length_in_scalar_cosine_similarity : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal data_a_in_scalar_cosine_similarity : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_b_in_scalar_cosine_similarity : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_scalar_cosine_similarity  : std_logic_vector(DATA_SIZE-1 downto 0);

  -- SCALAR EXPONENTIATOR
  -- CONTROL
  signal start_scalar_exponentiator : std_logic;
  signal ready_scalar_exponentiator : std_logic;

  -- DATA
  signal data_in_scalar_exponentiator  : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_scalar_exponentiator : std_logic_vector(DATA_SIZE-1 downto 0);

  -- SCALAR LOGARITHM
  -- CONTROL
  signal start_scalar_logarithm : std_logic;
  signal ready_scalar_logarithm : std_logic;

  -- DATA
  signal data_in_scalar_logarithm  : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_scalar_logarithm : std_logic_vector(DATA_SIZE-1 downto 0);

  -- SCALAR LOGISTIC
  -- CONTROL
  signal start_scalar_logistic : std_logic;
  signal ready_scalar_logistic : std_logic;

  -- DATA
  signal data_in_scalar_logistic  : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_scalar_logistic : std_logic_vector(DATA_SIZE-1 downto 0);

  -- CONTROL
  signal start_scalar_multiplication : std_logic;
  signal ready_scalar_multiplication : std_logic;

  signal data_in_enable_scalar_multiplication : std_logic;

  signal data_out_enable_scalar_multiplication : std_logic;

  -- DATA
  signal length_in_scalar_multiplication : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal data_in_scalar_multiplication   : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_scalar_multiplication  : std_logic_vector(DATA_SIZE-1 downto 0);

  -- SCALAR ONEPLUS
  -- CONTROL
  signal start_scalar_oneplus : std_logic;
  signal ready_scalar_oneplus : std_logic;

  -- DATA
  signal data_in_scalar_oneplus  : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_scalar_oneplus : std_logic_vector(DATA_SIZE-1 downto 0);

  -- SCALAR SINH
  -- CONTROL
  signal start_scalar_sinh : std_logic;
  signal ready_scalar_sinh : std_logic;

  -- DATA
  signal data_in_scalar_sinh  : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_scalar_sinh : std_logic_vector(DATA_SIZE-1 downto 0);

  -- CONTROL
  signal start_scalar_softmax : std_logic;
  signal ready_scalar_softmax : std_logic;

  signal data_in_enable_scalar_softmax : std_logic;

  signal data_out_enable_scalar_softmax : std_logic;

  -- DATA
  signal length_in_scalar_softmax : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal data_in_scalar_softmax   : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_scalar_softmax  : std_logic_vector(DATA_SIZE-1 downto 0);

  -- CONTROL
  signal start_scalar_summation : std_logic;
  signal ready_scalar_summation : std_logic;

  signal data_in_enable_scalar_summation : std_logic;

  signal data_out_enable_scalar_summation : std_logic;

  -- DATA
  signal length_in_scalar_summation : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal data_in_scalar_summation   : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_scalar_summation  : std_logic_vector(DATA_SIZE-1 downto 0);

  -- SCALAR TANH
  -- CONTROL
  signal start_scalar_tanh : std_logic;
  signal ready_scalar_tanh : std_logic;

  -- DATA
  signal data_in_scalar_tanh  : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_scalar_tanh : std_logic_vector(DATA_SIZE-1 downto 0);

  -----------------------------------------------------------------------
  -- VECTOR
  -----------------------------------------------------------------------

  -- VECTOR COSH
  -- CONTROL
  signal start_vector_cosh : std_logic;
  signal ready_vector_cosh : std_logic;

  signal data_in_enable_vector_cosh : std_logic;

  signal data_out_enable_vector_cosh : std_logic;

  -- DATA
  signal size_in_vector_cosh  : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal data_in_vector_cosh  : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_vector_cosh : std_logic_vector(DATA_SIZE-1 downto 0);

  -- VECTOR EXPONENTIATOR
  -- CONTROL
  signal start_vector_exponentiator : std_logic;
  signal ready_vector_exponentiator : std_logic;

  signal data_in_enable_vector_exponentiator : std_logic;

  signal data_out_enable_vector_exponentiator : std_logic;

  -- DATA
  signal size_in_vector_exponentiator  : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal data_in_vector_exponentiator  : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_vector_exponentiator : std_logic_vector(DATA_SIZE-1 downto 0);

  -- VECTOR LOGARITHM
  -- CONTROL
  signal start_vector_logarithm : std_logic;
  signal ready_vector_logarithm : std_logic;

  signal data_in_enable_vector_logarithm : std_logic;

  signal data_out_enable_vector_logarithm : std_logic;

  -- DATA
  signal size_in_vector_logarithm  : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal data_in_vector_logarithm  : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_vector_logarithm : std_logic_vector(DATA_SIZE-1 downto 0);

  -- VECTOR LOGISTIC
  -- CONTROL
  signal start_vector_logistic : std_logic;
  signal ready_vector_logistic : std_logic;

  signal data_in_enable_vector_logistic : std_logic;

  signal data_out_enable_vector_logistic : std_logic;

  -- DATA
  signal size_in_vector_logistic  : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal data_in_vector_logistic  : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_vector_logistic : std_logic_vector(DATA_SIZE-1 downto 0);

  -- VECTOR ONEPLUS
  -- CONTROL
  signal start_vector_oneplus : std_logic;
  signal ready_vector_oneplus : std_logic;

  signal data_in_enable_vector_oneplus : std_logic;

  signal data_out_enable_vector_oneplus : std_logic;

  -- DATA
  signal size_in_vector_oneplus  : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal data_in_vector_oneplus  : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_vector_oneplus : std_logic_vector(DATA_SIZE-1 downto 0);

  -- VECTOR SINH
  -- CONTROL
  signal start_vector_sinh : std_logic;
  signal ready_vector_sinh : std_logic;

  signal data_in_enable_vector_sinh : std_logic;

  signal data_out_enable_vector_sinh : std_logic;

  -- DATA
  signal size_in_vector_sinh  : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal data_in_vector_sinh  : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_vector_sinh : std_logic_vector(DATA_SIZE-1 downto 0);

  -- VECTOR TANH
  -- CONTROL
  signal start_vector_tanh : std_logic;
  signal ready_vector_tanh : std_logic;

  signal data_in_enable_vector_tanh : std_logic;

  signal data_out_enable_vector_tanh : std_logic;

  -- DATA
  signal size_in_vector_tanh  : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal data_in_vector_tanh  : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_vector_tanh : std_logic_vector(DATA_SIZE-1 downto 0);

  -----------------------------------------------------------------------
  -- MATRIX
  -----------------------------------------------------------------------

  -- MATRIX COSH
  -- CONTROL
  signal start_matrix_cosh : std_logic;
  signal ready_matrix_cosh : std_logic;

  signal data_in_i_enable_matrix_cosh : std_logic;
  signal data_in_j_enable_matrix_cosh : std_logic;

  signal data_out_i_enable_matrix_cosh : std_logic;
  signal data_out_j_enable_matrix_cosh : std_logic;

  -- DATA
  signal size_i_in_matrix_cosh : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal size_j_in_matrix_cosh : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal data_in_matrix_cosh   : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_matrix_cosh  : std_logic_vector(DATA_SIZE-1 downto 0);

  -- MATRIX EXPONENTIATOR
  -- CONTROL
  signal start_matrix_exponentiator : std_logic;
  signal ready_matrix_exponentiator : std_logic;

  signal data_in_i_enable_matrix_exponentiator : std_logic;
  signal data_in_j_enable_matrix_exponentiator : std_logic;

  signal data_out_i_enable_matrix_exponentiator : std_logic;
  signal data_out_j_enable_matrix_exponentiator : std_logic;

  -- DATA
  signal size_i_in_matrix_exponentiator : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal size_j_in_matrix_exponentiator : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal data_in_matrix_exponentiator   : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_matrix_exponentiator  : std_logic_vector(DATA_SIZE-1 downto 0);

  -- MATRIX LOGARITHM
  -- CONTROL
  signal start_matrix_logarithm : std_logic;
  signal ready_matrix_logarithm : std_logic;

  signal data_in_i_enable_matrix_logarithm : std_logic;
  signal data_in_j_enable_matrix_logarithm : std_logic;

  signal data_out_i_enable_matrix_logarithm : std_logic;
  signal data_out_j_enable_matrix_logarithm : std_logic;

  -- DATA
  signal size_i_in_matrix_logarithm : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal size_j_in_matrix_logarithm : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal data_in_matrix_logarithm   : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_matrix_logarithm  : std_logic_vector(DATA_SIZE-1 downto 0);

  -- MATRIX LOGISTIC
  -- CONTROL
  signal start_matrix_logistic : std_logic;
  signal ready_matrix_logistic : std_logic;

  signal data_in_i_enable_matrix_logistic : std_logic;
  signal data_in_j_enable_matrix_logistic : std_logic;

  signal data_out_i_enable_matrix_logistic : std_logic;
  signal data_out_j_enable_matrix_logistic : std_logic;

  -- DATA
  signal size_i_in_matrix_logistic : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal size_j_in_matrix_logistic : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal data_in_matrix_logistic   : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_matrix_logistic  : std_logic_vector(DATA_SIZE-1 downto 0);

  -- MATRIX ONEPLUS
  -- CONTROL
  signal start_matrix_oneplus : std_logic;
  signal ready_matrix_oneplus : std_logic;

  signal data_in_i_enable_matrix_oneplus : std_logic;
  signal data_in_j_enable_matrix_oneplus : std_logic;

  signal data_out_i_enable_matrix_oneplus : std_logic;
  signal data_out_j_enable_matrix_oneplus : std_logic;

  -- DATA
  signal size_i_in_matrix_oneplus : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal size_j_in_matrix_oneplus : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal data_in_matrix_oneplus   : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_matrix_oneplus  : std_logic_vector(DATA_SIZE-1 downto 0);

  -- MATRIX SINH
  -- CONTROL
  signal start_matrix_sinh : std_logic;
  signal ready_matrix_sinh : std_logic;

  signal data_in_i_enable_matrix_sinh : std_logic;
  signal data_in_j_enable_matrix_sinh : std_logic;

  signal data_out_i_enable_matrix_sinh : std_logic;
  signal data_out_j_enable_matrix_sinh : std_logic;

  -- DATA
  signal size_i_in_matrix_sinh : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal size_j_in_matrix_sinh : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal data_in_matrix_sinh   : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_matrix_sinh  : std_logic_vector(DATA_SIZE-1 downto 0);

  -- MATRIX TANH
  -- CONTROL
  signal start_matrix_tanh : std_logic;
  signal ready_matrix_tanh : std_logic;

  signal data_in_i_enable_matrix_tanh : std_logic;
  signal data_in_j_enable_matrix_tanh : std_logic;

  signal data_out_i_enable_matrix_tanh : std_logic;
  signal data_out_j_enable_matrix_tanh : std_logic;

  -- DATA
  signal size_i_in_matrix_tanh : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal size_j_in_matrix_tanh : std_logic_vector(CONTROL_SIZE-1 downto 0);
  signal data_in_matrix_tanh   : std_logic_vector(DATA_SIZE-1 downto 0);
  signal data_out_matrix_tanh  : std_logic_vector(DATA_SIZE-1 downto 0);

begin

  -----------------------------------------------------------------------
  -- Body
  -----------------------------------------------------------------------

  function_stimulus : ntm_function_stimulus
    generic map (
      -- SYSTEM-SIZE
      DATA_SIZE    => DATA_SIZE,
      CONTROL_SIZE => CONTROL_SIZE,

      X => X,
      Y => Y,
      N => N,
      W => W,
      L => L,
      R => R
      )
    port map (
      -- GLOBAL
      CLK => CLK,
      RST => RST,

      -----------------------------------------------------------------------
      -- STIMULUS SCALAR
      -----------------------------------------------------------------------

      -- SCALAR COSH
      -- CONTROL
      SCALAR_COSH_START => start_scalar_cosh,
      SCALAR_COSH_READY => ready_scalar_cosh,

      -- DATA
      SCALAR_COSH_DATA_IN  => data_in_scalar_cosh,
      SCALAR_COSH_DATA_OUT => data_out_scalar_cosh,

      -- SCALAR EXPONENTIATOR
      -- CONTROL
      SCALAR_EXPONENTIATOR_START => start_scalar_exponentiator,
      SCALAR_EXPONENTIATOR_READY => ready_scalar_exponentiator,

      -- DATA
      SCALAR_EXPONENTIATOR_DATA_IN  => data_in_scalar_exponentiator,
      SCALAR_EXPONENTIATOR_DATA_OUT => data_out_scalar_exponentiator,

      -- SCALAR LOGARITHM
      -- CONTROL
      SCALAR_LOGARITHM_START => start_scalar_logarithm,
      SCALAR_LOGARITHM_READY => ready_scalar_logarithm,

      -- DATA
      SCALAR_LOGARITHM_DATA_IN  => data_in_scalar_logarithm,
      SCALAR_LOGARITHM_DATA_OUT => data_out_scalar_logarithm,

      -- SCALAR LOGISTIC
      -- CONTROL
      SCALAR_LOGISTIC_START => start_scalar_logistic,
      SCALAR_LOGISTIC_READY => ready_scalar_logistic,

      -- DATA
      SCALAR_LOGISTIC_DATA_IN  => data_in_scalar_logistic,
      SCALAR_LOGISTIC_DATA_OUT => data_out_scalar_logistic,

      -- SCALAR ONEPLUS
      -- CONTROL
      SCALAR_ONEPLUS_START => start_scalar_oneplus,
      SCALAR_ONEPLUS_READY => ready_scalar_oneplus,

      -- DATA
      SCALAR_ONEPLUS_DATA_IN  => data_in_scalar_oneplus,
      SCALAR_ONEPLUS_DATA_OUT => data_out_scalar_oneplus,

      -- SCALAR SINH
      -- CONTROL
      SCALAR_SINH_START => start_scalar_sinh,
      SCALAR_SINH_READY => ready_scalar_sinh,

      -- DATA
      SCALAR_SINH_DATA_IN  => data_in_scalar_sinh,
      SCALAR_SINH_DATA_OUT => data_out_scalar_sinh,

      -- SCALAR TANH
      -- CONTROL
      SCALAR_TANH_START => start_scalar_tanh,
      SCALAR_TANH_READY => ready_scalar_tanh,

      -- DATA
      SCALAR_TANH_DATA_IN  => data_in_scalar_tanh,
      SCALAR_TANH_DATA_OUT => data_out_scalar_tanh,

      -----------------------------------------------------------------------
      -- STIMULUS VECTOR
      -----------------------------------------------------------------------

      -- VECTOR COSH
      -- CONTROL
      VECTOR_COSH_START => start_vector_cosh,
      VECTOR_COSH_READY => ready_vector_cosh,

      VECTOR_COSH_DATA_IN_ENABLE => data_in_enable_vector_cosh,

      VECTOR_COSH_DATA_OUT_ENABLE => data_out_enable_vector_cosh,

      -- DATA
      VECTOR_COSH_SIZE_IN  => size_in_vector_cosh,
      VECTOR_COSH_DATA_IN  => data_in_vector_cosh,
      VECTOR_COSH_DATA_OUT => data_out_vector_cosh,

      -- VECTOR EXPONENTIATOR
      -- CONTROL
      VECTOR_EXPONENTIATOR_START => start_vector_exponentiator,
      VECTOR_EXPONENTIATOR_READY => ready_vector_exponentiator,

      VECTOR_EXPONENTIATOR_DATA_IN_ENABLE => data_in_enable_vector_exponentiator,

      VECTOR_EXPONENTIATOR_DATA_OUT_ENABLE => data_out_enable_vector_exponentiator,

      -- DATA
      VECTOR_EXPONENTIATOR_SIZE_IN  => size_in_vector_exponentiator,
      VECTOR_EXPONENTIATOR_DATA_IN  => data_in_vector_exponentiator,
      VECTOR_EXPONENTIATOR_DATA_OUT => data_out_vector_exponentiator,

      -- VECTOR LOGARITHM
      -- CONTROL
      VECTOR_LOGARITHM_START => start_vector_logarithm,
      VECTOR_LOGARITHM_READY => ready_vector_logarithm,

      VECTOR_LOGARITHM_DATA_IN_ENABLE => data_in_enable_vector_logarithm,

      VECTOR_LOGARITHM_DATA_OUT_ENABLE => data_out_enable_vector_logarithm,

      -- DATA
      VECTOR_LOGARITHM_SIZE_IN  => size_in_vector_logarithm,
      VECTOR_LOGARITHM_DATA_IN  => data_in_vector_logarithm,
      VECTOR_LOGARITHM_DATA_OUT => data_out_vector_logarithm,

      -- VECTOR LOGISTIC
      -- CONTROL
      VECTOR_LOGISTIC_START => start_vector_logistic,
      VECTOR_LOGISTIC_READY => ready_vector_logistic,

      VECTOR_LOGISTIC_DATA_IN_ENABLE => data_in_enable_vector_logistic,

      VECTOR_LOGISTIC_DATA_OUT_ENABLE => data_out_enable_vector_logistic,

      -- DATA
      VECTOR_LOGISTIC_SIZE_IN  => size_in_vector_logistic,
      VECTOR_LOGISTIC_DATA_IN  => data_in_vector_logistic,
      VECTOR_LOGISTIC_DATA_OUT => data_out_vector_logistic,

      -- VECTOR ONEPLUS
      -- CONTROL
      VECTOR_ONEPLUS_START => start_vector_oneplus,
      VECTOR_ONEPLUS_READY => ready_vector_oneplus,

      VECTOR_ONEPLUS_DATA_IN_ENABLE => data_in_enable_vector_oneplus,

      VECTOR_ONEPLUS_DATA_OUT_ENABLE => data_out_enable_vector_oneplus,

      -- DATA
      VECTOR_ONEPLUS_SIZE_IN  => size_in_vector_oneplus,
      VECTOR_ONEPLUS_DATA_IN  => data_in_vector_oneplus,
      VECTOR_ONEPLUS_DATA_OUT => data_out_vector_oneplus,

      -- VECTOR SINH
      -- CONTROL
      VECTOR_SINH_START => start_vector_sinh,
      VECTOR_SINH_READY => ready_vector_sinh,

      VECTOR_SINH_DATA_IN_ENABLE => data_in_enable_vector_sinh,

      VECTOR_SINH_DATA_OUT_ENABLE => data_out_enable_vector_sinh,

      -- DATA
      VECTOR_SINH_SIZE_IN  => size_in_vector_sinh,
      VECTOR_SINH_DATA_IN  => data_in_vector_sinh,
      VECTOR_SINH_DATA_OUT => data_out_vector_sinh,

      -- VECTOR TANH
      -- CONTROL
      VECTOR_TANH_START => start_vector_tanh,
      VECTOR_TANH_READY => ready_vector_tanh,

      VECTOR_TANH_DATA_IN_ENABLE => data_in_enable_vector_tanh,

      VECTOR_TANH_DATA_OUT_ENABLE => data_out_enable_vector_tanh,

      -- DATA
      VECTOR_TANH_SIZE_IN  => size_in_vector_tanh,
      VECTOR_TANH_DATA_IN  => data_in_vector_tanh,
      VECTOR_TANH_DATA_OUT => data_out_vector_tanh,

      -----------------------------------------------------------------------
      -- STIMULUS MATRIX
      -----------------------------------------------------------------------

      -- MATRIX COSH
      -- CONTROL
      MATRIX_COSH_START => start_matrix_cosh,
      MATRIX_COSH_READY => ready_matrix_cosh,

      MATRIX_COSH_DATA_IN_I_ENABLE => data_in_i_enable_matrix_cosh,
      MATRIX_COSH_DATA_IN_J_ENABLE => data_in_j_enable_matrix_cosh,

      MATRIX_COSH_DATA_OUT_I_ENABLE => data_out_i_enable_matrix_cosh,
      MATRIX_COSH_DATA_OUT_J_ENABLE => data_out_j_enable_matrix_cosh,

      -- DATA
      MATRIX_COSH_SIZE_I_IN => size_i_in_matrix_cosh,
      MATRIX_COSH_SIZE_J_IN => size_j_in_matrix_cosh,
      MATRIX_COSH_DATA_IN   => data_in_matrix_cosh,
      MATRIX_COSH_DATA_OUT  => data_out_matrix_cosh,

      -- MATRIX EXPONENTIATOR
      -- CONTROL
      MATRIX_EXPONENTIATOR_START => start_matrix_exponentiator,
      MATRIX_EXPONENTIATOR_READY => ready_matrix_exponentiator,

      MATRIX_EXPONENTIATOR_DATA_IN_I_ENABLE => data_in_i_enable_matrix_exponentiator,
      MATRIX_EXPONENTIATOR_DATA_IN_J_ENABLE => data_in_j_enable_matrix_exponentiator,

      MATRIX_EXPONENTIATOR_DATA_OUT_I_ENABLE => data_out_i_enable_matrix_exponentiator,
      MATRIX_EXPONENTIATOR_DATA_OUT_J_ENABLE => data_out_j_enable_matrix_exponentiator,

      -- DATA
      MATRIX_EXPONENTIATOR_SIZE_I_IN => size_i_in_matrix_exponentiator,
      MATRIX_EXPONENTIATOR_SIZE_J_IN => size_j_in_matrix_exponentiator,
      MATRIX_EXPONENTIATOR_DATA_IN   => data_in_matrix_exponentiator,
      MATRIX_EXPONENTIATOR_DATA_OUT  => data_out_matrix_exponentiator,

      -- MATRIX LOGARITHM
      -- CONTROL
      MATRIX_LOGARITHM_START => start_matrix_logarithm,
      MATRIX_LOGARITHM_READY => ready_matrix_logarithm,

      MATRIX_LOGARITHM_DATA_IN_I_ENABLE => data_in_i_enable_matrix_logarithm,
      MATRIX_LOGARITHM_DATA_IN_J_ENABLE => data_in_j_enable_matrix_logarithm,

      MATRIX_LOGARITHM_DATA_OUT_I_ENABLE => data_out_i_enable_matrix_logarithm,
      MATRIX_LOGARITHM_DATA_OUT_J_ENABLE => data_out_j_enable_matrix_logarithm,

      -- DATA
      MATRIX_LOGARITHM_SIZE_I_IN => size_i_in_matrix_logarithm,
      MATRIX_LOGARITHM_SIZE_J_IN => size_j_in_matrix_logarithm,
      MATRIX_LOGARITHM_DATA_IN   => data_in_matrix_logarithm,
      MATRIX_LOGARITHM_DATA_OUT  => data_out_matrix_logarithm,

      -- MATRIX LOGISTIC
      -- CONTROL
      MATRIX_LOGISTIC_START => start_matrix_logistic,
      MATRIX_LOGISTIC_READY => ready_matrix_logistic,

      MATRIX_LOGISTIC_DATA_IN_I_ENABLE => data_in_i_enable_matrix_logistic,
      MATRIX_LOGISTIC_DATA_IN_J_ENABLE => data_in_j_enable_matrix_logistic,

      MATRIX_LOGISTIC_DATA_OUT_I_ENABLE => data_out_i_enable_matrix_logistic,
      MATRIX_LOGISTIC_DATA_OUT_J_ENABLE => data_out_j_enable_matrix_logistic,

      -- DATA
      MATRIX_LOGISTIC_SIZE_I_IN => size_i_in_matrix_logistic,
      MATRIX_LOGISTIC_SIZE_J_IN => size_j_in_matrix_logistic,
      MATRIX_LOGISTIC_DATA_IN   => data_in_matrix_logistic,
      MATRIX_LOGISTIC_DATA_OUT  => data_out_matrix_logistic,

      -- MATRIX ONEPLUS
      -- CONTROL
      MATRIX_ONEPLUS_START => start_matrix_oneplus,
      MATRIX_ONEPLUS_READY => ready_matrix_oneplus,

      MATRIX_ONEPLUS_DATA_IN_I_ENABLE => data_in_i_enable_matrix_oneplus,
      MATRIX_ONEPLUS_DATA_IN_J_ENABLE => data_in_j_enable_matrix_oneplus,

      MATRIX_ONEPLUS_DATA_OUT_I_ENABLE => data_out_i_enable_matrix_oneplus,
      MATRIX_ONEPLUS_DATA_OUT_J_ENABLE => data_out_j_enable_matrix_oneplus,

      -- DATA
      MATRIX_ONEPLUS_SIZE_I_IN => size_i_in_matrix_oneplus,
      MATRIX_ONEPLUS_SIZE_J_IN => size_j_in_matrix_oneplus,
      MATRIX_ONEPLUS_DATA_IN   => data_in_matrix_oneplus,
      MATRIX_ONEPLUS_DATA_OUT  => data_out_matrix_oneplus,

      -- MATRIX SINH
      -- CONTROL
      MATRIX_SINH_START => start_matrix_sinh,
      MATRIX_SINH_READY => ready_matrix_sinh,

      MATRIX_SINH_DATA_IN_I_ENABLE => data_in_i_enable_matrix_sinh,
      MATRIX_SINH_DATA_IN_J_ENABLE => data_in_j_enable_matrix_sinh,

      MATRIX_SINH_DATA_OUT_I_ENABLE => data_out_i_enable_matrix_sinh,
      MATRIX_SINH_DATA_OUT_J_ENABLE => data_out_j_enable_matrix_sinh,

      -- DATA
      MATRIX_SINH_SIZE_I_IN => size_i_in_matrix_sinh,
      MATRIX_SINH_SIZE_J_IN => size_j_in_matrix_sinh,
      MATRIX_SINH_DATA_IN   => data_in_matrix_sinh,
      MATRIX_SINH_DATA_OUT  => data_out_matrix_sinh,

      -- MATRIX TANH
      -- CONTROL
      MATRIX_TANH_START => start_matrix_tanh,
      MATRIX_TANH_READY => ready_matrix_tanh,

      MATRIX_TANH_DATA_IN_I_ENABLE => data_in_i_enable_matrix_tanh,
      MATRIX_TANH_DATA_IN_J_ENABLE => data_in_j_enable_matrix_tanh,

      MATRIX_TANH_DATA_OUT_I_ENABLE => data_out_i_enable_matrix_tanh,
      MATRIX_TANH_DATA_OUT_J_ENABLE => data_out_j_enable_matrix_tanh,

      -- DATA
      MATRIX_TANH_SIZE_I_IN => size_i_in_matrix_tanh,
      MATRIX_TANH_SIZE_J_IN => size_j_in_matrix_tanh,
      MATRIX_TANH_DATA_IN   => data_in_matrix_tanh,
      MATRIX_TANH_DATA_OUT  => data_out_matrix_tanh
      );

  -----------------------------------------------------------------------
  -- SCALAR
  -----------------------------------------------------------------------

  -- SCALAR COSH
  ntm_scalar_cosh_function_test : if (ENABLE_NTM_SCALAR_COSH_TEST) generate
    scalar_cosh_function : ntm_scalar_cosh_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_scalar_cosh,
        READY => ready_scalar_cosh,

        -- DATA
        DATA_IN  => data_in_scalar_cosh,
        DATA_OUT => data_out_scalar_cosh
        );
  end generate ntm_scalar_cosh_function_test;

  -- SCALAR EXPONENTIATOR
  ntm_scalar_exponentiator_function_test : if (ENABLE_NTM_SCALAR_EXPONENTIATOR_TEST) generate
    scalar_exponentiator_function : ntm_scalar_exponentiator_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_scalar_exponentiator,
        READY => ready_scalar_exponentiator,

        -- DATA
        DATA_IN  => data_in_scalar_exponentiator,
        DATA_OUT => data_out_scalar_exponentiator
        );
  end generate ntm_scalar_exponentiator_function_test;

  -- SCALAR LOGARITHM
  ntm_scalar_logarithm_function_test : if (ENABLE_NTM_SCALAR_LOGARITHM_TEST) generate
    scalar_logarithm_function : ntm_scalar_logarithm_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_scalar_logarithm,
        READY => ready_scalar_logarithm,

        -- DATA
        DATA_IN  => data_in_scalar_logarithm,
        DATA_OUT => data_out_scalar_logarithm
        );
  end generate ntm_scalar_logarithm_function_test;

  -- SCALAR LOGISTIC
  ntm_scalar_logistic_function_test : if (ENABLE_NTM_SCALAR_LOGISTIC_TEST) generate
    scalar_logistic_function : ntm_scalar_logistic_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_scalar_logistic,
        READY => ready_scalar_logistic,

        -- DATA
        DATA_IN  => data_in_scalar_logistic,
        DATA_OUT => data_out_scalar_logistic
        );
  end generate ntm_scalar_logistic_function_test;

  -- SCALAR ONEPLUS
  ntm_scalar_oneplus_function_test : if (ENABLE_NTM_SCALAR_ONEPLUS_TEST) generate
    scalar_oneplus_function : ntm_scalar_oneplus_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_scalar_oneplus,
        READY => ready_scalar_oneplus,

        -- DATA
        DATA_IN  => data_in_scalar_oneplus,
        DATA_OUT => data_out_scalar_oneplus
        );
  end generate ntm_scalar_oneplus_function_test;

  -- SCALAR SINH
  ntm_scalar_sinh_function_test : if (ENABLE_NTM_SCALAR_SINH_TEST) generate
    scalar_sinh_function : ntm_scalar_sinh_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_scalar_sinh,
        READY => ready_scalar_sinh,

        -- DATA
        DATA_IN  => data_in_scalar_sinh,
        DATA_OUT => data_out_scalar_sinh
        );
  end generate ntm_scalar_sinh_function_test;

  -- SCALAR TANH
  ntm_scalar_tanh_function_test : if (ENABLE_NTM_SCALAR_TANH_TEST) generate
    scalar_tanh_function : ntm_scalar_tanh_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_scalar_tanh,
        READY => ready_scalar_tanh,

        -- DATA
        DATA_IN  => data_in_scalar_tanh,
        DATA_OUT => data_out_scalar_tanh
        );
  end generate ntm_scalar_tanh_function_test;

  -----------------------------------------------------------------------
  -- VECTOR
  -----------------------------------------------------------------------

  -- VECTOR COSH
  ntm_vector_cosh_function_test : if (ENABLE_NTM_VECTOR_COSH_TEST) generate
    vector_cosh_function : ntm_vector_cosh_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_vector_cosh,
        READY => ready_vector_cosh,

        DATA_IN_ENABLE => data_in_enable_vector_cosh,

        DATA_OUT_ENABLE => data_out_enable_vector_cosh,

        -- DATA
        SIZE_IN  => size_in_vector_cosh,
        DATA_IN  => data_in_vector_cosh,
        DATA_OUT => data_out_vector_cosh
        );
  end generate ntm_vector_cosh_function_test;

  -- VECTOR EXPONENTIATOR
  ntm_vector_exponentiator_function_test : if (ENABLE_NTM_VECTOR_EXPONENTIATOR_TEST) generate
    vector_exponentiator_function : ntm_vector_exponentiator_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_vector_exponentiator,
        READY => ready_vector_exponentiator,

        DATA_IN_ENABLE => data_in_enable_vector_exponentiator,

        DATA_OUT_ENABLE => data_out_enable_vector_exponentiator,

        -- DATA
        SIZE_IN  => size_in_vector_exponentiator,
        DATA_IN  => data_in_vector_exponentiator,
        DATA_OUT => data_out_vector_exponentiator
        );
  end generate ntm_vector_exponentiator_function_test;

  -- VECTOR LOGARITHM
  ntm_vector_logarithm_function_test : if (ENABLE_NTM_VECTOR_LOGARITHM_TEST) generate
    vector_logarithm_function : ntm_vector_logarithm_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_vector_logarithm,
        READY => ready_vector_logarithm,

        DATA_IN_ENABLE => data_in_enable_vector_logarithm,

        DATA_OUT_ENABLE => data_out_enable_vector_logarithm,

        -- DATA
        SIZE_IN  => size_in_vector_logarithm,
        DATA_IN  => data_in_vector_logarithm,
        DATA_OUT => data_out_vector_logarithm
        );
  end generate ntm_vector_logarithm_function_test;

  -- VECTOR LOGISTIC
  ntm_vector_logistic_function_test : if (ENABLE_NTM_VECTOR_LOGISTIC_TEST) generate
    vector_logistic_function : ntm_vector_logistic_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_vector_logistic,
        READY => ready_vector_logistic,

        DATA_IN_ENABLE => data_in_enable_vector_logistic,

        DATA_OUT_ENABLE => data_out_enable_vector_logistic,

        -- DATA
        SIZE_IN  => size_in_vector_logistic,
        DATA_IN  => data_in_vector_logistic,
        DATA_OUT => data_out_vector_logistic
        );
  end generate ntm_vector_logistic_function_test;

  -- VECTOR ONEPLUS
  ntm_vector_oneplus_function_test : if (ENABLE_NTM_VECTOR_ONEPLUS_TEST) generate
    vector_oneplus_function : ntm_vector_oneplus_function
      generic map (

        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_vector_oneplus,
        READY => ready_vector_oneplus,

        DATA_IN_ENABLE => data_in_enable_vector_oneplus,

        DATA_OUT_ENABLE => data_out_enable_vector_oneplus,

        -- DATA
        SIZE_IN  => size_in_vector_oneplus,
        DATA_IN  => data_in_vector_oneplus,
        DATA_OUT => data_out_vector_oneplus
        );
  end generate ntm_vector_oneplus_function_test;

  -- VECTOR SINH
  ntm_vector_sinh_function_test : if (ENABLE_NTM_VECTOR_SINH_TEST) generate
    vector_sinh_function : ntm_vector_sinh_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_vector_sinh,
        READY => ready_vector_sinh,

        DATA_IN_ENABLE => data_in_enable_vector_sinh,

        DATA_OUT_ENABLE => data_out_enable_vector_sinh,

        -- DATA
        SIZE_IN  => size_in_vector_sinh,
        DATA_IN  => data_in_vector_sinh,
        DATA_OUT => data_out_vector_sinh
        );
  end generate ntm_vector_sinh_function_test;

  -- VECTOR TANH
  ntm_vector_tanh_function_test : if (ENABLE_NTM_VECTOR_TANH_TEST) generate
    vector_tanh_function : ntm_vector_tanh_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_vector_tanh,
        READY => ready_vector_tanh,

        DATA_IN_ENABLE => data_in_enable_vector_tanh,

        DATA_OUT_ENABLE => data_out_enable_vector_tanh,

        -- DATA
        SIZE_IN  => size_in_vector_tanh,
        DATA_IN  => data_in_vector_tanh,
        DATA_OUT => data_out_vector_tanh
        );
  end generate ntm_vector_tanh_function_test;

  -----------------------------------------------------------------------
  -- MATRIX
  -----------------------------------------------------------------------

  -- MATRIX COSH
  ntm_matrix_cosh_function_test : if (ENABLE_NTM_MATRIX_COSH_TEST) generate
    matrix_cosh_function : ntm_matrix_cosh_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_matrix_cosh,
        READY => ready_matrix_cosh,

        DATA_IN_I_ENABLE => data_in_i_enable_matrix_cosh,
        DATA_IN_J_ENABLE => data_in_j_enable_matrix_cosh,

        DATA_OUT_I_ENABLE => data_out_i_enable_matrix_cosh,
        DATA_OUT_J_ENABLE => data_out_j_enable_matrix_cosh,

        -- DATA
        SIZE_I_IN => size_i_in_matrix_cosh,
        SIZE_J_IN => size_j_in_matrix_cosh,
        DATA_IN   => data_in_matrix_cosh,
        DATA_OUT  => data_out_matrix_cosh
        );
  end generate ntm_matrix_cosh_function_test;

  -- MATRIX EXPONENTIATOR
  ntm_matrix_exponentiator_function_test : if (ENABLE_NTM_MATRIX_EXPONENTIATOR_TEST) generate
    matrix_exponentiator_function : ntm_matrix_exponentiator_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_matrix_exponentiator,
        READY => ready_matrix_exponentiator,

        DATA_IN_I_ENABLE => data_in_i_enable_matrix_exponentiator,
        DATA_IN_J_ENABLE => data_in_j_enable_matrix_exponentiator,

        DATA_OUT_I_ENABLE => data_out_i_enable_matrix_exponentiator,
        DATA_OUT_J_ENABLE => data_out_j_enable_matrix_exponentiator,

        -- DATA
        SIZE_I_IN => size_i_in_matrix_exponentiator,
        SIZE_J_IN => size_j_in_matrix_exponentiator,
        DATA_IN   => data_in_matrix_exponentiator,
        DATA_OUT  => data_out_matrix_exponentiator
        );
  end generate ntm_matrix_exponentiator_function_test;

  -- MATRIX LOGARITHM
  ntm_matrix_logarithm_function_test : if (ENABLE_NTM_MATRIX_LOGARITHM_TEST) generate
    matrix_logarithm_function : ntm_matrix_logarithm_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_matrix_logarithm,
        READY => ready_matrix_logarithm,

        DATA_IN_I_ENABLE => data_in_i_enable_matrix_logarithm,
        DATA_IN_J_ENABLE => data_in_j_enable_matrix_logarithm,

        DATA_OUT_I_ENABLE => data_out_i_enable_matrix_logarithm,
        DATA_OUT_J_ENABLE => data_out_j_enable_matrix_logarithm,

        -- DATA
        SIZE_I_IN => size_i_in_matrix_logarithm,
        SIZE_J_IN => size_j_in_matrix_logarithm,
        DATA_IN   => data_in_matrix_logarithm,
        DATA_OUT  => data_out_matrix_logarithm
        );
  end generate ntm_matrix_logarithm_function_test;

  -- MATRIX LOGISTIC
  ntm_matrix_logistic_function_test : if (ENABLE_NTM_MATRIX_LOGISTIC_TEST) generate
    matrix_logistic_function : ntm_matrix_logistic_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_matrix_logistic,
        READY => ready_matrix_logistic,

        DATA_IN_I_ENABLE => data_in_i_enable_matrix_logistic,
        DATA_IN_J_ENABLE => data_in_j_enable_matrix_logistic,

        DATA_OUT_I_ENABLE => data_out_i_enable_matrix_logistic,
        DATA_OUT_J_ENABLE => data_out_j_enable_matrix_logistic,

        -- DATA
        SIZE_I_IN => size_i_in_matrix_logistic,
        SIZE_J_IN => size_j_in_matrix_logistic,
        DATA_IN   => data_in_matrix_logistic,
        DATA_OUT  => data_out_matrix_logistic
        );
  end generate ntm_matrix_logistic_function_test;

  -- MATRIX ONEPLUS
  ntm_matrix_oneplus_function_test : if (ENABLE_NTM_MATRIX_ONEPLUS_TEST) generate
    matrix_oneplus_function : ntm_matrix_oneplus_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_matrix_oneplus,
        READY => ready_matrix_oneplus,

        DATA_IN_I_ENABLE => data_in_i_enable_matrix_oneplus,
        DATA_IN_J_ENABLE => data_in_j_enable_matrix_oneplus,

        DATA_OUT_I_ENABLE => data_out_i_enable_matrix_oneplus,
        DATA_OUT_J_ENABLE => data_out_j_enable_matrix_oneplus,

        -- DATA
        SIZE_I_IN => size_i_in_matrix_oneplus,
        SIZE_J_IN => size_j_in_matrix_oneplus,
        DATA_IN   => data_in_matrix_oneplus,
        DATA_OUT  => data_out_matrix_oneplus
        );
  end generate ntm_matrix_oneplus_function_test;

  -- MATRIX SINH
  ntm_matrix_sinh_function_test : if (ENABLE_NTM_MATRIX_SINH_TEST) generate
    matrix_sinh_function : ntm_matrix_sinh_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_matrix_sinh,
        READY => ready_matrix_sinh,

        DATA_IN_I_ENABLE => data_in_i_enable_matrix_sinh,
        DATA_IN_J_ENABLE => data_in_j_enable_matrix_sinh,

        DATA_OUT_I_ENABLE => data_out_i_enable_matrix_sinh,
        DATA_OUT_J_ENABLE => data_out_j_enable_matrix_sinh,

        -- DATA
        SIZE_I_IN => size_i_in_matrix_sinh,
        SIZE_J_IN => size_j_in_matrix_sinh,
        DATA_IN   => data_in_matrix_sinh,
        DATA_OUT  => data_out_matrix_sinh
        );
  end generate ntm_matrix_sinh_function_test;

  -- MATRIX TANH
  ntm_matrix_tanh_function_test : if (ENABLE_NTM_MATRIX_TANH_TEST) generate
    matrix_tanh_function : ntm_matrix_tanh_function
      generic map (
        DATA_SIZE    => DATA_SIZE,
        CONTROL_SIZE => CONTROL_SIZE
        )
      port map (
        -- GLOBAL
        CLK => CLK,
        RST => RST,

        -- CONTROL
        START => start_matrix_tanh,
        READY => ready_matrix_tanh,

        DATA_IN_I_ENABLE => data_in_i_enable_matrix_tanh,
        DATA_IN_J_ENABLE => data_in_j_enable_matrix_tanh,

        DATA_OUT_I_ENABLE => data_out_i_enable_matrix_tanh,
        DATA_OUT_J_ENABLE => data_out_j_enable_matrix_tanh,

        -- DATA
        SIZE_I_IN => size_i_in_matrix_tanh,
        SIZE_J_IN => size_j_in_matrix_tanh,
        DATA_IN   => data_in_matrix_tanh,
        DATA_OUT  => data_out_matrix_tanh
        );
  end generate ntm_matrix_tanh_function_test;

end ntm_function_testbench_architecture;
