--------------------------------------------------------------------------------
--                                            __ _      _     _               --
--                                           / _(_)    | |   | |              --
--                __ _ _   _  ___  ___ _ __ | |_ _  ___| | __| |              --
--               / _` | | | |/ _ \/ _ \ '_ \|  _| |/ _ \ |/ _` |              --
--              | (_| | |_| |  __/  __/ | | | | | |  __/ | (_| |              --
--               \__, |\__,_|\___|\___|_| |_|_| |_|\___|_|\__,_|              --
--                  | |                                                       --
--                  |_|                                                       --
--                                                                            --
--                                                                            --
--              Peripheral-NTM for MPSoC                                      --
--              Neural Turing Machine for MPSoC                               --
--                                                                            --
--------------------------------------------------------------------------------

-- Copyright (c) 2020-2021 by the author(s)
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
-- THE SOFTWARE.
--
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.ntm_math_pkg.all;

package ntm_core_pkg is

  -----------------------------------------------------------------------
  -- Constants
  -----------------------------------------------------------------------

  -----------------------------------------------------------------------
  -- Components
  -----------------------------------------------------------------------

  -----------------------------------------------------------------------
  -- READ HEADS
  -----------------------------------------------------------------------

  component ntm_reading is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      M_IN_ENABLE  : in  std_logic;
      R_OUT_ENABLE : out std_logic;

      -- DATA
      W_IN  : in  std_logic_vector(DATA_SIZE-1 downto 0);
      M_IN  : in  std_logic_vector(DATA_SIZE-1 downto 0);
      R_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  -----------------------------------------------------------------------
  -- WRITE HEADS
  -----------------------------------------------------------------------

  component ntm_writing is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      M_IN_ENABLE  : in std_logic;
      A_IN_ENABLE  : in std_logic;
      M_OUT_ENABLE : in std_logic;

      -- DATA
      M_IN  : in std_logic_vector(DATA_SIZE-1 downto 0);
      A_IN  : in std_logic_vector(DATA_SIZE-1 downto 0);
      W_IN  : in std_logic_vector(DATA_SIZE-1 downto 0);
      M_OUT : in std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component ntm_erasing is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      M_IN_ENABLE  : in std_logic;
      E_IN_ENABLE  : in std_logic;
      M_OUT_ENABLE : in std_logic;

      -- DATA
      M_IN  : in std_logic_vector(DATA_SIZE-1 downto 0);
      E_IN  : in std_logic_vector(DATA_SIZE-1 downto 0);
      W_IN  : in std_logic_vector(DATA_SIZE-1 downto 0);
      M_OUT : in std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  -----------------------------------------------------------------------
  -- MEMORY
  -----------------------------------------------------------------------

  component ntm_content_based_addressing is
    generic (
      I : integer := 64;
      J : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      K_IN_ENABLE : in std_logic; -- for j in 0 to J-1

      M_IN_I_ENABLE : in std_logic; -- for i in 0 to I-1
      M_IN_J_ENABLE : in std_logic; -- for j in 0 to J-1

      C_OUT_ENABLE : out std_logic; -- for i in 0 to I-1

      -- DATA
      K_IN    : in std_logic_vector(DATA_SIZE-1 downto 0);
      M_IN    : in std_logic_vector(DATA_SIZE-1 downto 0);
      BETA_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      C_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component ntm_addressing is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      K_IN_ENABLE : in std_logic; -- for k in 0 to W-1
      S_IN_ENABLE : in std_logic; -- for k in 0 to W-1

      M_IN_J_ENABLE : in std_logic; -- for j in 0 to N-1
      M_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1

      W_IN_ENABLE  : in  std_logic; -- for j in 0 to N-1
      W_OUT_ENABLE : out std_logic; -- for j in 0 to N-1

      -- DATA
      K_IN     : in std_logic_vector(DATA_SIZE-1 downto 0);
      BETA_IN  : in std_logic_vector(DATA_SIZE-1 downto 0);
      G_IN     : in std_logic_vector(DATA_SIZE-1 downto 0);
      S_IN     : in std_logic_vector(DATA_SIZE-1 downto 0);
      GAMMA_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      M_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      W_IN  : in  std_logic_vector(DATA_SIZE-1 downto 0);
      W_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  -----------------------------------------------------------------------
  -- TOP
  -----------------------------------------------------------------------

  component ntm_top is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      X_IN_ENABLE : in std_logic; -- for x in 0 to X-1

      Y_OUT_ENABLE : out std_logic; -- for y in 0 to Y-1

      -- DATA
      X_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      Y_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component ntm_interface_vector is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      -- Key Vector
      WK_IN_L_ENABLE : in std_logic; -- for l in 0 to L-1
      WK_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1

      K_OUT_ENABLE : out std_logic; -- for k in 0 to W-1

      -- Key Strength
      WBETA_IN_ENABLE : in std_logic; -- for l in 0 to L-1

      -- Interpolation Gate
      WG_IN_ENABLE : in std_logic; -- for l in 0 to L-1

      -- Shift Weighting
      WS_IN_L_ENABLE : in std_logic; -- for l in 0 to L-1
      WS_IN_J_ENABLE : in std_logic; -- for j in 0 to N-1

      S_OUT_ENABLE : out std_logic; -- for j in 0 to N-1

      -- Sharpening
      WGAMMA_IN_ENABLE : in std_logic; -- for l in 0 to L-1

      -- Hidden State
      H_IN_ENABLE : in std_logic; -- for l in 0 to L-1

      -- DATA
      WK_IN     : in std_logic_vector(DATA_SIZE-1 downto 0);
      WBETA_IN  : in std_logic_vector(DATA_SIZE-1 downto 0);
      WG_IN     : in std_logic_vector(DATA_SIZE-1 downto 0);
      WS_IN     : in std_logic_vector(DATA_SIZE-1 downto 0);
      WGAMMA_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      H_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      K_OUT     : out std_logic_vector(DATA_SIZE-1 downto 0);
      BETA_OUT  : out std_logic_vector(DATA_SIZE-1 downto 0);
      G_OUT     : out std_logic_vector(DATA_SIZE-1 downto 0);
      S_OUT     : out std_logic_vector(DATA_SIZE-1 downto 0);
      GAMMA_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component ntm_output_vector is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      K_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1
      K_IN_Y_ENABLE : in std_logic; -- for y in 0 to Y-1
      K_IN_K_ENABLE : in std_logic; -- for k in 0 to W-1

      R_IN_I_ENABLE : in std_logic; -- for i in 0 to R-1
      R_IN_K_ENABLE : in std_logic; -- for j in 0 to W-1

      NU_IN_ENABLE : in std_logic; -- for y in 0 to Y-1

      Y_OUT_ENABLE : in std_logic; -- for y in 0 to Y-1

      -- DATA
      K_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      R_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      NU_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      Y_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

  component ntm_controller_output_vector is
    generic (
      X : integer := 64;
      Y : integer := 64;
      N : integer := 64;
      W : integer := 64;
      L : integer := 64;

      DATA_SIZE : integer := 512
    );
    port (
      -- GLOBAL
      CLK : in std_logic;
      RST : in std_logic;

      -- CONTROL
      START : in  std_logic;
      READY : out std_logic;

      U_IN_Y_ENABLE : in std_logic; -- for y in 0 to Y-1
      U_IN_L_ENABLE : in std_logic; -- for l in 0 to L-1

      H_IN_ENABLE : in std_logic; -- for l in 0 to L-1

      NU_ENABLE_OUT : out std_logic; -- for j in 0 to Y-1

      -- DATA
      U_IN : in std_logic_vector(DATA_SIZE-1 downto 0);
      H_IN : in std_logic_vector(DATA_SIZE-1 downto 0);

      NU_OUT : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
  end component;

end ntm_core_pkg;
